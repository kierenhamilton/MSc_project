module DEC (
  input [31:0] PC,
  input [31:0] rs1,
  input [31:0] rs2,
  );

  endmodule
