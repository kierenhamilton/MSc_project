module branLog ();
endmodule
