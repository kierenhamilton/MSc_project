module progMem ();
endmodule
