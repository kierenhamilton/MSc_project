module progCounter();
endmodule
