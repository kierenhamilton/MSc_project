module ram ();
endmodule
