module regMem ();
endmodule
